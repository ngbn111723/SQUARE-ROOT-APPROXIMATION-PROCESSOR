library verilog;
use verilog.vl_types.all;
entity ADD_SUB_module_vlg_vec_tst is
end ADD_SUB_module_vlg_vec_tst;
