library verilog;
use verilog.vl_types.all;
entity AU_vlg_vec_tst is
end AU_vlg_vec_tst;
