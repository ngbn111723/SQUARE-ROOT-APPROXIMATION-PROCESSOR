library verilog;
use verilog.vl_types.all;
entity AU_1_vlg_vec_tst is
end AU_1_vlg_vec_tst;
