library verilog;
use verilog.vl_types.all;
entity Datapath_pipelining_vlg_vec_tst is
end Datapath_pipelining_vlg_vec_tst;
