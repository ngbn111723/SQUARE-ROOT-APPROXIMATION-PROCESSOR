library verilog;
use verilog.vl_types.all;
entity AU_2_vlg_vec_tst is
end AU_2_vlg_vec_tst;
